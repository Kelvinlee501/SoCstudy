NORMAL_TEST
