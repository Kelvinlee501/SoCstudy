
`define P_CLK_PERIOD   10
`define PARAM_TEMPLETE 0
