
`define VIP_ADDR_WIDTH 32
`define VIP_DATA_WIDTH 32
