////////////////////////////////////
//
//
//
////////////////////////////////////

module src_templete #(
	parameter			PARAM = 1	
) (
	input						I_CLK,
	input						I_RESETn
);

endmodule
