
	// Design Parameter
	parameter		P_CLOCK_PERIOD		= 10;
	parameter		PARAM_TEMPLETE		= 0;

	// Verification Parameter - Don't change

	// Monitor Control Parameter

	// VIP Control Parameter

	// test Control Parameter
