
	initial begin
		warning_count = 0;
		error_count = 0;
	end

