
//=========================================================
// apb4 Master
//=========================================================
//
// VIP interface
	assign apb4_m_vip.pclk    = top.clk;
	assign apb4_m_vip.presetn = top.resetn;

	//please describe VIP interface
	
//=========================================================
// AXI4 Slave
//=========================================================


//=========================================================
// I2C
//=========================================================
