

module apb4_m_monitor;


endmodule
