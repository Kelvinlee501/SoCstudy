

module axi_s_monitor;


endmodule
