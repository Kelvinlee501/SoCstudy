	integer			local_error_cnt;
