
	integer	warning_count;
	integer error_count;
